/*Input Interface*/

`ifndef INPINF
 `define INPINF
 `include "primitives.vh"

module inpinf #(parameter XB = 10,
				parameter YB = 10,
				parameter PB = 8)
	(/*AUTOARG*/
	// Outputs
	px_in_ready, col_count, row_count,
	// Inputs
	clk, rst, cfg_width, cfg_height, px_in_data, px_in_valid
	);

	//Globals
	input clk;
	input rst;

	//Frame Config
	input [XB-1:0] cfg_width;
	input [YB-1:0] cfg_height;
	
	//Input Data
	input [PB-1:0] px_in_data;
	input 		   px_in_valid; 

	output 		   px_in_ready;
	output [XB-1:0] col_count;
	output [YB-1:0] row_count;
	
	

	
	//Input fifo to collect pixels
	//Inputs to Fifo
	wire 		   inq_wr, inq_rd;
	wire [PB-1:0]  inq_datain;

	//Outputs
	wire 		   inq_full, inq_al_full;
	wire 		   inq_emty, inq_al_emty;
	wire [PB-1:0]  inq_dataout;
	
	
	
	hw_fifo inp_fifo (
					  // Outputs
					  .wr_full			(inq_full),
					  .wr_almost_full	(inq_al_full),
					  .rd_data			(inq_dataout),
					  .rd_empty			(inq_emty),
					  .rd_almost_empty	(inq_al_emty),
					  // Inputs
					  .clk				(clk),
					  .rst				(rst),
					  .wr_push			(inq_wr),
					  .wr_data			(inq_datain),
					  .rd_pop			(inq_rd));
	
	//Loading data into input Fifo
	assign px_in_ready = ~inq_full;	
	assign inq_wr = px_in_valid & px_in_ready;
	assign inq_datain = px_in_data;
	assign inq_rd = 1'b1;
	
	//Column Count - Counts number of pixels coming in
	reg [XB-1:0]   col_count;
	wire 		   inc_col_count;
	wire 		   rst_col_count;
	
	assign inc_col_count = inq_rd;
	assign rst_col_count = (col_count >= cfg_width) || rst;
	`EN_ASYNC_RST_MSFF(col_count, col_count+1'b1, clk, inc_col_count, rst_col_count)

	//Row Count - Counts number of rows
	reg [YB-1:0]   row_count;
	wire 		   inc_row_count;
	wire 		   rst_row_count;
	assign inc_row_count = (col_count == cfg_width);
	assign rst_row_count = (row_count >= cfg_height) || rst;
	`EN_ASYNC_RST_MSFF(row_count, row_count+1'b1, clk, inc_row_count, rst_row_count)

	
endmodule // inpInf
`endif


   
	
